`include "test_package.sv"

module tb_int_cpu_jump ();
  import test_package :: *;

  logic clk, reset, uart_rx, uart_tx;
  test_clock test_clock(clk);
  assign uart_rx = 1'b1; // no signal

  mother_board #(.WAIT(8), .FILENAME("")) mother_board(.*);

  function automatic void init_mem_restart_cpu(input [31:0] init_vals[]);
    int n = init_vals.size();
    mother_board.rom.mem = '{default: '{default: '0}};
    for (int i = 0; i < n; i++) mother_board.rom.mem[i] = init_vals[i];

    reset = 1'b1;
    #RESET_PERIOD;
    reset = 1'b0;
    #(PERIOD_PER_INSTRUCT*n);
  endfunction

  logic [15:0][31:0] x;
  assign x = mother_board.cpu.gr_file.x;

  initial begin
    // ----------------------------------------------------------------------------------------------------
    // jalr
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___1___4___0___2 // jalr ---- x[4] = pc + 1; pc = x[1]
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd7, x[1]); // jump addr
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump
    `check32(32'd4, x[4]); // back addr

    // ----------------------------------------------------------------------------------------------------
    // jeq
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h001___0___0___4___0___0 // addi ---- x[4] = x[0] + 1
      , 32'h000___4___1___0___0___3 // jeq  ---- if (x[4] == 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___0___4___0___0 // addi ---- x[4] = x[0] + 0
      , 32'h000___4___1___0___0___3 // jeq  ---- if (x[4] == 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'hFFF___0___0___4___0___0 // addi ---- x[4] = x[0] + (-1)
      , 32'h000___4___1___0___0___3 // jeq  ---- if (x[4] == 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    // ----------------------------------------------------------------------------------------------------
    // jneq
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h001___0___0___4___0___0 // addi ---- x[4] = x[0] + 1
      , 32'h000___4___1___0___1___3 // jneq ---- if (x[4] != 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___0___4___0___0 // addi ---- x[4] = x[0] + 0
      , 32'h000___4___1___0___1___3 // jneq ---- if (x[4] != 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'hFFF___0___0___4___0___0 // addi ---- x[4] = x[0] + (-1)
      , 32'h000___4___1___0___1___3 // jneq ---- if (x[4] != 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    // ----------------------------------------------------------------------------------------------------
    // jge
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h001___0___0___4___0___0 // addi ---- x[4] = x[0] + 1
      , 32'h000___4___1___0___2___3 // jneq ---- if (x[4] >= 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___0___4___0___0 // addi ---- x[4] = x[0] + 0
      , 32'h000___4___1___0___2___3 // jneq ---- if (x[4] >= 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'hFFF___0___0___4___0___0 // addi ---- x[4] = x[0] + (-1)
      , 32'h000___4___1___0___2___3 // jneq ---- if (x[4] >= 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    // ----------------------------------------------------------------------------------------------------
    // jlt
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h001___0___0___4___0___0 // addi ---- x[4] = x[0] + 1
      , 32'h000___4___1___0___3___3 // jneq ---- if (x[4] < 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___0___4___0___0 // addi ---- x[4] = x[0] + 0
      , 32'h000___4___1___0___3___3 // jneq ---- if (x[4] < 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'hFFF___0___0___4___0___0 // addi ---- x[4] = x[0] + (-1)
      , 32'h000___4___1___0___3___3 // jneq ---- if (x[4] < 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump


    // ----------------------------------------------------------------------------------------------------
    // jgt
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h001___0___0___4___0___0 // addi ---- x[4] = x[0] + 1
      , 32'h000___4___1___0___4___3 // jneq ---- if (x[4] > 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___0___4___0___0 // addi ---- x[4] = x[0] + 0
      , 32'h000___4___1___0___4___3 // jneq ---- if (x[4] > 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'hFFF___0___0___4___0___0 // addi ---- x[4] = x[0] + (-1)
      , 32'h000___4___1___0___4___3 // jneq ---- if (x[4] > 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump


    // ----------------------------------------------------------------------------------------------------
    // jle
    // ----------------------------------------------------------------------------------------------------

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h001___0___0___4___0___0 // addi ---- x[4] = x[0] + 1
      , 32'h000___4___1___0___5___3 // jneq ---- if (x[4] <= 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd1, x[2]); // is not jump
    `check32(32'd0, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'h000___0___0___4___0___0 // addi ---- x[4] = x[0] + 0
      , 32'h000___4___1___0___5___3 // jneq ---- if (x[4] <= 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump

    init_mem_restart_cpu('{
        //  imm  rs2 rs1 rd  opt opcode
        32'h007___0___0___1___0___0 // addi ---- x[1] = x[0] + 7
      , 32'h000___0___0___2___0___0 // addi ---- x[2] = x[0] + 0
      , 32'h000___0___0___3___0___0 // addi ---- x[3] = x[0] + 0
      , 32'hFFF___0___0___4___0___0 // addi ---- x[4] = x[0] + (-1)
      , 32'h000___4___1___0___5___3 // jneq ---- if (x[4] <= 0) {pc = x[1]}
      , 32'h001___0___0___2___0___0 // addi ---- x[2] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
      , 32'h001___0___0___3___0___0 // addi ---- x[3] = x[0] + 1
      , 32'h000___0___0___0___0___A // halt
    });
    `check32(32'd0, x[2]); // is not jump
    `check32(32'd1, x[3]); // is jump
  end
endmodule
